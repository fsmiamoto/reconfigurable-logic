lpm_counter1_inst : lpm_counter1 PORT MAP (
		aclr	 => aclr_sig,
		clock	 => clock_sig,
		q	 => q_sig
	);
