-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Full Version
-- Created on Fri Mar 26 17:31:33 2021

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY LineFollower IS
    PORT (
        clock : IN STD_LOGIC;
        reset : IN STD_LOGIC := '0';
        left_sensor : IN STD_LOGIC := '0';
        right_sensor : IN STD_LOGIC := '0';
        left_motor_1 : OUT STD_LOGIC;
        left_motor_2 : OUT STD_LOGIC;
        right_motor_1 : OUT STD_LOGIC;
        right_motor_2 : OUT STD_LOGIC
    );
END LineFollower;

ARCHITECTURE BEHAVIOR OF LineFollower IS
    TYPE type_fstate IS (Stopped,Turning_Right,Turning_Left,Forward);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
    SIGNAL reg_left_motor_1 : STD_LOGIC := '0';
    SIGNAL reg_left_motor_2 : STD_LOGIC := '0';
    SIGNAL reg_right_motor_1 : STD_LOGIC := '0';
    SIGNAL reg_right_motor_2 : STD_LOGIC := '0';
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,left_sensor,right_sensor,reg_left_motor_1,reg_left_motor_2,reg_right_motor_1,reg_right_motor_2)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= Forward;
            reg_left_motor_1 <= '0';
            reg_left_motor_2 <= '0';
            reg_right_motor_1 <= '0';
            reg_right_motor_2 <= '0';
            left_motor_1 <= '0';
            left_motor_2 <= '0';
            right_motor_1 <= '0';
            right_motor_2 <= '0';
        ELSE
            reg_left_motor_1 <= '0';
            reg_left_motor_2 <= '0';
            reg_right_motor_1 <= '0';
            reg_right_motor_2 <= '0';
            left_motor_1 <= '0';
            left_motor_2 <= '0';
            right_motor_1 <= '0';
            right_motor_2 <= '0';
            CASE fstate IS
                WHEN Stopped =>
                    IF (((left_sensor = '1') AND (right_sensor = '1'))) THEN
                        reg_fstate <= Forward;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Stopped;
                    END IF;

                    reg_right_motor_1 <= '0';

                    reg_left_motor_1 <= '0';

                    reg_right_motor_2 <= '0';

                    reg_left_motor_2 <= '0';
                WHEN Turning_Right =>
                    IF ((NOT((left_sensor = '1')) AND NOT((right_sensor = '1')))) THEN
                        reg_fstate <= Stopped;
                    ELSIF (((left_sensor = '1') AND (right_sensor = '1'))) THEN
                        reg_fstate <= Forward;
                    ELSIF ((NOT((left_sensor = '1')) AND (right_sensor = '1'))) THEN
                        reg_fstate <= Turning_Left;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Turning_Right;
                    END IF;

                    reg_right_motor_1 <= '0';

                    reg_left_motor_1 <= '1';

                    reg_right_motor_2 <= '0';

                    reg_left_motor_2 <= '0';
                WHEN Turning_Left =>
                    IF ((NOT((left_sensor = '1')) AND NOT((right_sensor = '1')))) THEN
                        reg_fstate <= Stopped;
                    ELSIF (((left_sensor = '1') AND NOT((right_sensor = '1')))) THEN
                        reg_fstate <= Turning_Right;
                    ELSIF (((left_sensor = '1') AND (right_sensor = '1'))) THEN
                        reg_fstate <= Forward;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Turning_Left;
                    END IF;

                    reg_right_motor_1 <= '1';

                    reg_left_motor_1 <= '0';

                    reg_right_motor_2 <= '0';

                    reg_left_motor_2 <= '0';
                WHEN Forward =>
                    IF (((left_sensor = '1') AND NOT((right_sensor = '1')))) THEN
                        reg_fstate <= Turning_Right;
                    ELSIF ((NOT((left_sensor = '1')) AND NOT((right_sensor = '1')))) THEN
                        reg_fstate <= Stopped;
                    ELSIF ((NOT((left_sensor = '1')) AND (right_sensor = '1'))) THEN
                        reg_fstate <= Turning_Left;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Forward;
                    END IF;

                    reg_right_motor_1 <= '1';

                    reg_left_motor_1 <= '1';

                    reg_right_motor_2 <= '1';

                    reg_left_motor_2 <= '1';
                WHEN OTHERS => 
                    reg_left_motor_1 <= 'X';
                    reg_left_motor_2 <= 'X';
                    reg_right_motor_1 <= 'X';
                    reg_right_motor_2 <= 'X';
                    report "Reach undefined state";
            END CASE;
            left_motor_1 <= reg_left_motor_1;
            left_motor_2 <= reg_left_motor_2;
            right_motor_1 <= reg_right_motor_1;
            right_motor_2 <= reg_right_motor_2;
        END IF;
    END PROCESS;
END BEHAVIOR;
