-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.


-- Generated by Quartus II 64-Bit Version 13.0 (Build Build 232 06/12/2013)
-- Created on Tue Mar 09 17:19:59 2021

StateMachine StateMachine_inst
(
	.clock(clock_sig) ,	// input  clock_sig
	.reset(reset_sig) ,	// input  reset_sig
	.direction(direction_sig) ,	// input  direction_sig
	.enable(enable_sig) ,	// input  enable_sig
	.output_1(output_1_sig) ,	// output  output_1_sig
	.output_2(output_2_sig) 	// output  output_2_sig
);

