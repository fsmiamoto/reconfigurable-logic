library verilog;
use verilog.vl_types.all;
entity RootMeanSquare_vlg_vec_tst is
end RootMeanSquare_vlg_vec_tst;
