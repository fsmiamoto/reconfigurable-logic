lpm_mult0_inst : lpm_mult0 PORT MAP (
		dataa	 => dataa_sig,
		result	 => result_sig
	);
