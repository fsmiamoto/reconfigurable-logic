lpm_counter0_inst : lpm_counter0 PORT MAP (
		clock	 => clock_sig,
		q	 => q_sig
	);
